`timescale 1ns / 1ps

module mixcolumnd(a,mcl);
input [127:0] a;
output [127:0] mcl;

wire [127:0] lut14,lut13,lut11,lut9;

     gm_lut14 q0( .a(a[127:120]),.c(lut14[127:120]) );
     gm_lut14 q1( .a(a[119:112]),.c(lut14[119:112]) );
     gm_lut14 q2( .a(a[111:104]),.c(lut14[111:104]) );
     gm_lut14 q3( .a(a[103:96]),.c(lut14[103:96]) );    
     gm_lut14 q4( .a(a[95:88]),.c(lut14[95:88]) );
     gm_lut14 q5( .a(a[87:80]),.c(lut14[87:80]) );
     gm_lut14 q6( .a(a[79:72]),.c(lut14[79:72]) );
     gm_lut14 q7( .a(a[71:64]),.c(lut14[71:64]) );     
     gm_lut14 q8( .a(a[63:56]),.c(lut14[63:56]) );
     gm_lut14 q9( .a(a[55:48]),.c(lut14[55:48]) );
     gm_lut14 q10(.a(a[47:40]),.c(lut14[47:40]) );
     gm_lut14 q11(.a(a[39:32]),.c(lut14[39:32]) );     
     gm_lut14 q12(.a(a[31:24]),.c(lut14[31:24]) );
     gm_lut14 q13(.a(a[23:16]),.c(lut14[23:16]) );
     gm_lut14 q14(.a(a[15:8]),.c(lut14[15:8]) );
     gm_lut14 q16(.a(a[7:0]),.c(lut14[7:0]) );

     gm_lut13 p0( .a(a[127:120]),.c(lut13[127:120]) );
     gm_lut13 p1( .a(a[119:112]),.c(lut13[119:112]) );
     gm_lut13 p2( .a(a[111:104]),.c(lut13[111:104]) );
     gm_lut13 p3( .a(a[103:96]),.c(lut13[103:96]) );   
     gm_lut13 p4( .a(a[95:88]),.c(lut13[95:88]) );
     gm_lut13 p5( .a(a[87:80]),.c(lut13[87:80]) );
     gm_lut13 p6( .a(a[79:72]),.c(lut13[79:72]) );
     gm_lut13 p7( .a(a[71:64]),.c(lut13[71:64]) );
     gm_lut13 p8( .a(a[63:56]),.c(lut13[63:56]) );
     gm_lut13 p9( .a(a[55:48]),.c(lut13[55:48]) );
     gm_lut13 p10(.a(a[47:40]),.c(lut13[47:40]) );
     gm_lut13 p11(.a(a[39:32]),.c(lut13[39:32]) );
     gm_lut13 p12(.a(a[31:24]),.c(lut13[31:24]) );
     gm_lut13 p13(.a(a[23:16]),.c(lut13[23:16]) );
     gm_lut13 p14(.a(a[15:8]),.c(lut13[15:8]) );
     gm_lut13 p16(.a(a[7:0]),.c(lut13[7:0]) );
     
     gm_lut11 r0( .a(a[127:120]),.c(lut11[127:120]) );
     gm_lut11 r1( .a(a[119:112]),.c(lut11[119:112]) );
     gm_lut11 r2( .a(a[111:104]),.c(lut11[111:104]) );
     gm_lut11 r3( .a(a[103:96]),.c(lut11[103:96]) );     
     gm_lut11 r4( .a(a[95:88]),.c(lut11[95:88]) );
     gm_lut11 r5( .a(a[87:80]),.c(lut11[87:80]) );
     gm_lut11 r6( .a(a[79:72]),.c(lut11[79:72]) );
     gm_lut11 r7( .a(a[71:64]),.c(lut11[71:64]) );     
     gm_lut11 r8( .a(a[63:56]),.c(lut11[63:56]) );
     gm_lut11 r9( .a(a[55:48]),.c(lut11[55:48]) );
     gm_lut11 r10(.a(a[47:40]),.c(lut11[47:40]) );
     gm_lut11 r11(.a(a[39:32]),.c(lut11[39:32]) );     
     gm_lut11 r12(.a(a[31:24]),.c(lut11[31:24]) );
     gm_lut11 r13(.a(a[23:16]),.c(lut11[23:16]) );
     gm_lut11 r14(.a(a[15:8]),.c(lut11[15:8]) );
     gm_lut11 r16(.a(a[7:0]),.c(lut11[7:0]) );
     
     gm_lut9 s0( .a(a[127:120]),.c(lut9[127:120]) );
     gm_lut9 s1( .a(a[119:112]),.c(lut9[119:112]) );
     gm_lut9 s2( .a(a[111:104]),.c(lut9[111:104]) );
     gm_lut9 s3( .a(a[103:96]),.c(lut9[103:96]) );     
     gm_lut9 s4( .a(a[95:88]),.c(lut9[95:88]) );
     gm_lut9 s5( .a(a[87:80]),.c(lut9[87:80]) );
     gm_lut9 s6( .a(a[79:72]),.c(lut9[79:72]) );
     gm_lut9 s7( .a(a[71:64]),.c(lut9[71:64]) );     
     gm_lut9 s8( .a(a[63:56]),.c(lut9[63:56]) );
     gm_lut9 s9( .a(a[55:48]),.c(lut9[55:48]) );
     gm_lut9 s10(.a(a[47:40]),.c(lut9[47:40]) );
     gm_lut9 s11(.a(a[39:32]),.c(lut9[39:32]) );     
     gm_lut9 s12(.a(a[31:24]),.c(lut9[31:24]) );
     gm_lut9 s13(.a(a[23:16]),.c(lut9[23:16]) );
     gm_lut9 s14(.a(a[15:8]),.c(lut9[15:8]) );
     gm_lut9 s16(.a(a[7:0]),.c(lut9[7:0]) );

assign mcl[127:120]= lut14[127:120] ^ lut11[119:112] ^ lut13[111:104] ^ lut9[103:96];
assign mcl[119:112]= lut14[119:112] ^ lut11[111:104] ^ lut13[103:96] ^ lut9[127:120];
assign mcl[111:104]= lut14[111:104] ^ lut11[103:96] ^ lut13[127:120] ^ lut9[119:112];
assign mcl[103:96]= lut14[103:96] ^ lut11[127:120] ^ lut13[119:112] ^ lut9[111:104];

assign mcl[95:88]= lut14[95:88] ^ lut11[87:80] ^ lut13[79:72] ^ lut9[71:64];
assign mcl[87:80]= lut14[87:80] ^ lut11[79:72] ^ lut13[71:64] ^ lut9[95:88];
assign mcl[79:72]= lut14[79:72] ^ lut11[71:64] ^ lut13[95:88] ^ lut9[87:80];
assign mcl[71:64]= lut14[71:64] ^ lut11[95:88] ^ lut13[87:80] ^ lut9[79:72];

assign mcl[63:56]= lut14[63:56] ^ lut11[55:48] ^ lut13[47:40] ^ lut9[39:32];
assign mcl[55:48]= lut14[55:48] ^ lut11[47:40] ^ lut13[39:32] ^ lut9[63:56];
assign mcl[47:40]= lut14[47:40] ^ lut11[39:32] ^ lut13[63:56] ^ lut9[55:48];
assign mcl[39:32]= lut14[39:32] ^ lut11[63:56] ^ lut13[55:48] ^ lut9[47:40];

assign mcl[31:24]= lut14[31:24] ^ lut11[23:16] ^ lut13[15:8] ^ lut9[7:0];
assign mcl[23:16]= lut14[23:16] ^ lut11[15:8] ^ lut13[7:0] ^ lut9[31:24];
assign mcl[15:8]= lut14[15:8] ^ lut11[7:0] ^ lut13[31:24] ^ lut9[23:16];
assign mcl[7:0]= lut14[7:0] ^ lut11[31:24] ^ lut13[23:16] ^ lut9[15:8];


endmodule
